module exec #(parameter OPCODE_WIDTH    =  4,
                        PMEM_ADDR_WIDTH = 12,
                        PMEM_WORD_WIDTH = 16,
                        IALU_WORD_WIDTH = 16,
                        REG_IDX_WIDTH   =  4,
                        PC_WIDTH        = 12,
                        PC_INCREMENT    =  2)
             (
             input                         clock,
             input                         reset,
             input                         in_act_ialu_add,
             input                         in_act_incr_pc_is_res,
             input                         in_act_jump_to_ialu_res,
             input                         in_act_write_res_to_reg,
             input  [       PC_WIDTH-1:0]  in_pc,
             input  [  REG_IDX_WIDTH-1:0]  in_res_reg_idx,
             input  [IALU_WORD_WIDTH-1:0]  in_src1,
             input  [IALU_WORD_WIDTH-1:0]  in_src2,
             output                        out_act_write_res_to_reg,
             output                        out_flush,
             output [PMEM_ADDR_WIDTH-1:0]  out_new_pc,
             output [IALU_WORD_WIDTH-1:0]  out_res,
             output [  REG_IDX_WIDTH-1:0]  out_res_reg_idx,
             output                        out_set_pc
             );

    // Sampled inputs
    reg                       act_ialu_add_sampled;
    reg                       act_incr_pc_is_res_sampled;
    reg                       act_jump_to_ialu_res_sampled;
    reg [       PC_WIDTH-1:0] pc_sampled;
    reg [IALU_WORD_WIDTH-1:0] src1_sampled;
    reg [IALU_WORD_WIDTH-1:0] src2_sampled;
    
    // ALU regs
    reg [IALU_WORD_WIDTH-1:0] ialu_res;
    
    
    // Register: sample inputs
    always @(posedge clock or posedge reset)
    begin
        if (!reset) begin
            act_ialu_add_sampled         <= in_act_ialu_add;
            act_incr_pc_is_res_sampled   <= in_act_incr_pc_is_res;
            act_jump_to_ialu_res_sampled <= in_act_jump_to_ialu_res;
            pc_sampled                   <= in_pc;
            src1_sampled                 <= in_src1;
            src2_sampled                 <= in_src2;
        end
        else begin
            act_ialu_add_sampled         <= 0;
            act_incr_pc_is_res_sampled   <= 0;
            act_jump_to_ialu_res_sampled <= 0;
            pc_sampled                   <= 0;
            src1_sampled                 <= 0;
            src2_sampled                 <= 0;
        end
    end

    // Register: pass through
    always @(posedge clock or posedge reset) begin
        if (!reset) begin
            out_act_write_res_to_reg <= in_act_write_res_to_reg;
            out_res_reg_idx          <= in_res_reg_idx;
        end
        else begin
            out_act_write_res_to_reg <= 0;
            out_res_reg_idx          <= 0;
        end
    end

    // ALU
    always @(*)
    begin
        // Integer addition
        if (act_ialu_add_sampled) begin
            ialu_res = src1_sampled + src2_sampled;
        end
        
        // default: do nothing
        else begin
            ialu_res = 0;
        end
    end

    // JUMP / BRANCH
    always @(*)
    begin
        // Trigger jump after getting 2nd instruction word with immedate target address
        if (act_jump_to_ialu_res_sampled) begin
            out_flush  = 1;
            out_set_pc = 1;
            out_new_pc = out_res[PMEM_ADDR_WIDTH-1:0];
        end
        else begin
            out_flush  = 0;
            out_set_pc = 0;
            out_new_pc = 0;
        end
    end

    // Multiplexer: forward either IALU result or incremented PC to result lane
    always @(*)
    begin
        if (act_incr_pc_is_res_sampled) begin
             out_res[IALU_WORD_WIDTH-1:PC_WIDTH] = 0;
             out_res[       PC_WIDTH-1:       0] = pc_sampled + PC_INCREMENT;
        end
        else begin
             out_res = ialu_res;           
        end
    end

endmodule

